module main
import os
import cp
fn main() {
	cp.run_cp(os.args)
}
