module mvutil

struct MvCommand{
	
}
