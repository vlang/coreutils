module main
import os
import cp
fn main() {
<<<<<<< HEAD
	run_cp(os.args)
	// 
=======
	cp.run_cp(os.args)
>>>>>>> e94acd3 (Rearranged modules to make the main executable of module main)
}
