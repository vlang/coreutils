module main

fn test_1() {
	println(@METHOD)
	assert true
}