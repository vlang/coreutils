module main
import os
import rm

// import src.rm.rmutil
fn main() {
	rm.run_rm(os.args)
}
