module pwd

pub struct UserInfo {
pub:
	username string
	uid      int
	gid      int
}
