module main

import os
import src.cp

fn main() {
	cp.run_cp(os.args)
}
