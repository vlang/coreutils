module main

import os
import src.rm

fn main() {
	rm.run_rm(os.args)
}
