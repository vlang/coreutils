module mvutil

struct MvCommand {
}
