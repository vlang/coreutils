module main

import os
import rm

fn main() {
	rm.run_rm(os.args)
}
