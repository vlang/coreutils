module mvutil

struct MvCommand {
}

fn (m MvCommand) run() {
	println(name)
}
