module main

import os
import src.rm

// import src.rm.rmutil
fn main() {
	rm.run_rm(os.args)
}
