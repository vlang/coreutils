module main

import os
import src.cp

fn main() {
	run_cp(os.args)
	// 
}
