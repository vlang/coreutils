module main

fn test_stub() {
	assert true
}
