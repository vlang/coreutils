module pwd
