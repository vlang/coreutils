module main
import os
import mv

fn main() {
	mv.run_mv(os.args)
}
