module main

import os
import src.mv

fn main() {
	mv.run_mv(os.args)
}
