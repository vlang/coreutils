module main

import os
import rmutil

fn main() {
	rmutil.run_rm(os.args)
}
