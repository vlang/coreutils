module main

fn main() {
	exit(1)
}
