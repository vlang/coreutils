module main

fn main() {
	exit(0)
}

